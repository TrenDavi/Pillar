module write
(
   input wire clk,
   input wire reset
);

endmodule
