module decode
(
   input wire clk,
   input wire reset
);
// Decode logic

// Register Fetch

endmodule
